----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    05:33:54 05/20/2014 
-- Design Name: 
-- Module Name:    VGACounter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;


entity VGACounter is
    Port ( CLK : in  STD_LOGIC;  -- Se asume a 50 MHz
           RST : in  STD_LOGIC;
           PBTON : in  STD_LOGIC;
           HS : out  STD_LOGIC;
           VS : out  STD_LOGIC;
           RGB : out  STD_LOGIC_VECTOR (11 downto 0)
     );
			  	
end VGACounter;

architecture Behavioral of VGACounter is
	-- Declaramos componentes
	COMPONENT BIN2BCD_0a999
	PORT(
		BIN : IN std_logic_vector(9 downto 0);          
		BCD2 : OUT std_logic_vector(3 downto 0);
		BCD1 : OUT std_logic_vector(3 downto 0);
		BCD0 : OUT std_logic_vector(3 downto 0)
		);
	END COMPONENT;
	
	COMPONENT vga_ctrl_640x480_60Hz
	PORT(
		rst : IN std_logic;
		clk : IN std_logic; 
		rgb_in : IN std_logic_vector(11 downto 0);          
		HS : OUT std_logic;
		VS : OUT std_logic;
		hcount : OUT std_logic_vector(10 downto 0);
		vcount : OUT std_logic_vector(10 downto 0);
		rgb_out : OUT std_logic_vector(11 downto 0);
		blank : OUT std_logic
		);
	END COMPONENT;
	
	COMPONENT Display 
	GENERIC ( LW: INTEGER:=10;
				 DW: INTEGER:=50;
				 DL: INTEGER:=100;
				 POSX: INTEGER:= 0;
				 POSY: INTEGER:= 0
         	); 
   PORT (  HCOUNT : in  STD_LOGIC_VECTOR (10 downto 0);
           VCOUNT : in  STD_LOGIC_VECTOR (10 downto 0);
           VALUE : in  STD_LOGIC_VECTOR (3 downto 0);
           PAINT : out  STD_LOGIC);
	end COMPONENT;
	
	COMPONENT AlphaNumerico
	GENERIC ( LW: INTEGER:=10;
				 DW: INTEGER:=50;
				 DL: INTEGER:=100;
				 POSX: INTEGER:= 0;
				 POSY: INTEGER:= 0
         	); 
	PORT(
		ALPHANUM : IN std_logic_vector(6 downto 0);
		HCOUNT : IN std_logic_vector(10 downto 0);
		VCOUNT : IN std_logic_vector(10 downto 0);          
		PAINT : OUT std_logic
		);
	END COMPONENT;
	
	-- Declaramos segnales
	signal hcount : STD_LOGIC_VECTOR (10 downto 0);
	signal vcount : STD_LOGIC_VECTOR (10 downto 0);
    signal paint2 : STD_LOGIC;
    signal paint1 : STD_LOGIC;
    signal paint0 : STD_LOGIC;
    
	signal rgb_aux1 : STD_LOGIC_VECTOR (2 downto 0);
	signal rgb_aux2 : STD_LOGIC_VECTOR (11 downto 0);
	signal rgb_aux3 : STD_LOGIC_VECTOR (11 downto 0);
	
	signal conteo : std_logic_vector(9 downto 0);
	signal unidades : std_logic_vector(3 downto 0);
	signal decenas : std_logic_vector(3 downto 0);
	signal centenas : std_logic_vector(3 downto 0);
	
	signal CLK_1Hz : STD_LOGIC:='0';
	signal clk_interno : STD_LOGIC:='0';
    signal cnt_pixeles: integer := 0;


	
begin

	Inst_vga_ctrl_640x480_60Hz: vga_ctrl_640x480_60Hz PORT MAP(
		rst => RST,
		clk => clk,
		rgb_in => rgb_aux3,
		HS => HS,
		VS => VS,
		hcount => hcount,
		vcount => vcount,
		rgb_out => rgb_aux2,
		blank => open
	);

    pixel_clk_stimulus: process(clk)
	begin
		if (clk'event and clk = '1') then
			clk_interno <= NOT clk_interno;
		end if;
	end process;
    --
	--CLK_DIV_60HZ: process (CLK)
	--	variable cnt: integer:= 0;
    --begin  
	--   if (CLK'event and CLK = '1') then
	--	if 	cnt = 416666 then
	--		clk_interno <= '1';
	--	elsif cnt = 833333 then
	--		clk_interno <= '0';
	--		cnt := 0;			
	--	else 
	--		cnt := cnt + 1;
	--	end if;
    --        
    --   end if;
    --end process;
	
	-- *****************************************************************************************************************
	-- Se comenta para la prueba (es dificil ver el resultado del incremento del contador cada segundo por simulacion)
	--
	-- CLK_DIV_1HZ: process(clk_interno)
	-- begin
	-- 	 if(clk_interno'event and clk_interno='1') then
	--		 if (count_clk = 5000000) then
	--			 count_clk <= 0;
	--			 CLK_1Hz <= not CLK_1Hz;
	--       	 else
	--			 count_clk <= count_clk + 1;
	--	     end if;
	--    end if;
	-- end process;
	-- *****************************************************************************************************************
	
	-- DYSPLAY_CONT: process(CLK_1Hz,RST)
	-- clk interno es el reloj de 50 MHz
	DYSPLAY_CONT: process(clk_interno,RST)

	begin
		if (RST='1') then
			conteo <= (others=>'0');
		elsif (clk_interno'event and clk_interno='1') then	-- elsif (CLK_1Hz'event and CLK_1Hz='1') then
			if(PBTON='1') then                 
                if cnt_pixeles = 420000 then 
              		if (conteo=999) then
				    	conteo <= (others=>'0');
				    else
					    conteo <= conteo + 1;
                    end if;
                    cnt_pixeles <= 0;
                else
                    cnt_pixeles <= cnt_pixeles + 1;
				end if;              
			else
				conteo <= conteo;
			end if;
		end if;
	end process;
	
	BIN2BCD: BIN2BCD_0a999 PORT MAP(
		BIN => conteo,
		BCD2 => centenas,
		BCD1 => decenas,
		BCD0 => unidades
	);
	
	Display2: Display  
	GENERIC MAP (
		LW => 40,
		DW => 200,
		DL => 320,
		POSX => 100,
		POSY => 80)
	PORT MAP(
		HCOUNT => hcount,
		VCOUNT => vcount,
		VALUE => centenas,
		PAINT => paint2
	);
	
	Display1: Display  
	GENERIC MAP (
		LW => 10,
		DW => 50,
		DL => 80,
		POSX => 345,
		POSY => 320)
	PORT MAP(
		HCOUNT => hcount,
		VCOUNT => vcount,
		VALUE => decenas,
		PAINT => paint1
	);
	
	Display0: Display 
	GENERIC MAP (
		LW => 20,
		DW => 100,
		DL => 160,
		POSX => 440,
		POSY => 240)
	PORT MAP(
		HCOUNT => hcount,
		VCOUNT => vcount,
		VALUE => unidades,
		PAINT => paint0
	);

	rgb_aux1 <= "110" when paint2='1' else
	            "001" when paint1='1' else
				"100" when paint0='1' else
				"000";
	rgb_aux3 <= rgb_aux1(2)&rgb_aux1(2)&rgb_aux1(2)&rgb_aux1(2)&rgb_aux1(1)&rgb_aux1(1)&rgb_aux1(1)&rgb_aux1(1)&rgb_aux1(0)&rgb_aux1(0)&rgb_aux1(0)&rgb_aux1(0);

	RGB <= rgb_aux2;
	
end Behavioral;

